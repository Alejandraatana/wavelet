--Alejandra Rodriguez Sanchez Ing. en Computacion
library ieee;

use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity senal is
   port(
           add: in std_logic_vector(7 downto 0);
           dat:out std_logic_vector(15 downto 0)
       );
end entity senal;
architecture beh of senal is
type data is array (0 to 255) of std_logic_vector(15 downto 0);
signal dato: data:=
               (
                  0=>"0000000000000000",
                  1=>"0001111000110001",
                  2=>"0001110010100010",
                  3=>"0010011101011011",
                  4=>"0010101011110110",
                  5=>"0010110011101110",
                  6=>"0010111000000101",
                  7=>"0011000001111101",
                  8=>"0011000011110010",
                  9=>"0011011011110110",
                 10=>"0011010111011101",
                 11=>"0100011100001010",
                 12=>"0011100001000001",
                 13=>"0100000100110011",
                 14=>"0100000100001110",
                 15=>"0100010000010000",
                 16=>"0101001001110000",
                 17=>"0100001101001110",
                 18=>"0101000010110000",
                 19=>"0101010001010000",
                 20=>"0101001100110001",
                 21=>"0100111000010010",
                 22=>"0101000101001000",
                 23=>"0100101111111111",
                 24=>"0101110111011101",
                 25=>"0101001111001111",
                 26=>"0101001101100110",
                 27=>"0100110110001110",
                 28=>"0101101110110100",
                 29=>"0100101110010101",
                 30=>"0100001001100100",
                 31=>"0101000001000010",
                 32=>"0100001100100011",
                 33=>"0011110010111100", 
                 34=>"0010001111011011", 
                 35=>"0010000110001010", 
                 36=>"0001101110110111",
                 37=>"0010010111110110",
                 38=>"0001010000011100",
                 39=>"0000111111001111",
                 40=>"0000111100100001",
                 41=>"0001000100101110",
                 42=>"0000101110101101",
                 43=>"0000111100001000",
                 44=>"0000101101100100",
                 45=>"0000010001110110",
                 46=>"0000100101111011",
                 47=>"0000000011111010",
                 48=>"0000101110110011",
                 49=>"0000011101111110",
                 50=>"0001000011001001",
                 51=>"0000001001101001",
                 52=>"0000101010011011",
                 53=>"0000011001111110",
                 54=>"0000011001010101",
                 55=>"0000001111000000",
                 56=>"0000000111110100",
                 57=>"0000100001000010",
                 58=>"0000100100110010",
                 59=>"0000101101010100",
                 60=>"0001001100001110",
                 61=>"0010001100001100",
                 62=>"0010010011110100",
                 63=>"0010110000010011",
                 64=>"0011111100010011",
                 65=>"0100000011101001",
                 66=>"0100000110001010",
                 67=>"0100100100010111",
                 68=>"0101011000010100",
                 69=>"0110111100010000",
                 70=>"0111010000111100",
                 71=>"0110000101110000",
                 72=>"0110101000111111",
                 73=>"0110110001110000",
                 74=>"0111011111110010",
                 75=>"0111101110110111",
                 76=>"0111110110111001",
                 77=>"0111111000100010",
                 78=>"0111011100000110",
                 79=>"0111111101101000",
                 80=>"0111110101001011",
                 81=>"0111110111010010",
                 82=>"0111000010010110",
                 83=>"0111100001100111",
                 84=>"0111001111000000",
                 85=>"0111000111100101",
                 86=>"0111101101100001",
                 87=>"0101111001000101",
                 88=>"0101101011001101",
                 89=>"0101011111110100",
                 90=>"0100100001010001",
                 91=>"0100011110011010",
                 92=>"0011110001011010",
                 93=>"0011000110001101",
                 94=>"0010110010111011",
                 95=>"0010110000010000",
                 96=>"0010001110011100",
                 97=>"0001111100100111",
                 98=>"0010000001000111",
                 99=>"0010000000001011",
                100=>"0001001000100001",
                101=>"0001010001110000",
                102=>"0001011001011100",
                103=>"0001000011111011",
                104=>"0001000011011111",
                105=>"0000101111100101",
                106=>"0000010001001011",
                107=>"0000011111110011",
                108=>"0000100101101011",
                109=>"0000011010111111",
                110=>"0000001101010100",
                111=>"0000010001101110",
                112=>"0000001111000110",
                113=>"0000101100010110",
                114=>"0001011110010001",
                115=>"0000100100001111",
                116=>"0000110011011110",
                117=>"0000111000000011",
                118=>"0010001101110100",
                119=>"0001010001001010",
                120=>"0001101001000101",
                121=>"0001011110010000",
                122=>"0001100100101100",
                123=>"0010100000110101",
                124=>"0010010100100011",
                125=>"0010101010000001",
                126=>"0010101100011100",
                127=>"0011000111110101",
                128=>"0011001000001101",
                129=>"0011101000101101",
                130=>"0100000001010001",
                131=>"0011111111010000",
                132=>"0100000111010110",
                133=>"0100101100110001",
                134=>"0101101001010110",
                135=>"0101001111010101",
                136=>"0100100011100001",
                137=>"0100111111111010",
                138=>"0110000100100111",
                139=>"0100111001001110",
                140=>"0101100100110000",
                141=>"0101010010110001",
                142=>"0101010111011010",
                143=>"0101101000001101",
                144=>"0101000001011001",
                145=>"0110000011100001",
                146=>"0100101001100101",
                147=>"0100111001111100",
                148=>"0100110000001110",
                149=>"0100100000001110",
                150=>"0100100110100011",
                151=>"0100011100100010",
                152=>"0011101011100110",
                153=>"0011111110110101",
                154=>"0011101011001111",
                155=>"0011100001011011",
                156=>"0011101011100010",
                157=>"0010101000011000",
                158=>"0011011111101111",
                159=>"0011011101100111",
                160=>"0001111100110000",
                161=>"0010000010011000",
                162=>"0001101110011111",
                163=>"0010010111001011",
                164=>"0001011101100001",
                165=>"0000111001011111",
                166=>"0000100100010001",
                167=>"0001101001100101",
                168=>"0000110011011011",
                169=>"0001001110001011",
                170=>"0000010101111001",
                171=>"0000011010111100",
                172=>"0000011101000001",
                173=>"0000101000101101",
                174=>"0000001100100011",
                175=>"0000101010110110",
                176=>"0000101110011011",
                177=>"0000100100000010",
                178=>"0000111010001010",
                179=>"0000110100000100",
                180=>"0001000101001011",
                181=>"0001011010000010",
                182=>"0001010100000111",
                183=>"0001111000001100",
                184=>"0010000011110100",
                185=>"0011010101011100",
                186=>"0001111101010010",
                187=>"0010010001010111",
                188=>"0010100110000010",
                189=>"0011111100101011",
                190=>"0011011101010011",
                191=>"0100001100001001",
                192=>"0100101100001110",
                193=>"0101001010110011",
                194=>"0100001101111010",
                195=>"0101000010001000",
                196=>"0100011101101001",
                197=>"0101001010110011",
                198=>"0100011100101100",
                199=>"0100101101110011",
                200=>"0101100000011110",
                201=>"0101001110010001",
                202=>"0101011110011111",
                203=>"0100111011011010",
                204=>"0110000000101011",
                205=>"0101010111101101",
                206=>"0101110110000010",
                207=>"0100111000111101",
                208=>"0101000011010110",
                209=>"0101000010101000",
                210=>"0101001010110101",
                211=>"0100111110011001",
                212=>"0100101011001011",
                213=>"0100100010010010",
                214=>"0100000111000111",
                215=>"0011110101110111",
                216=>"0011111000100011",
                217=>"0100011010001011",
                218=>"0010111101001111",
                219=>"0010111110010010",
                220=>"0010101111000001",
                221=>"0010100101010001",
                222=>"0010101110011000",
                223=>"0010000100100101",
                224=>"0001101110011001",
                225=>"0001111010101100",
                226=>"0001011011101001",
                227=>"0001001011111000",
                228=>"0000111101110011",
                229=>"0001101010010011",
                230=>"0000110101110100",
                231=>"0000011001010000",
                232=>"0000001011001101",
                233=>"0000110000100001",
                234=>"0000001011000000",
                235=>"0000010111000001",
                236=>"0000011110011100",
                237=>"0001000110110110",
                238=>"0001011010101000",
                239=>"0000011011011101",
                240=>"0000010000001110",
                241=>"0000100110000011",
                242=>"0001001001000101",
                243=>"0001111111011011",
                244=>"0001101011010110",
                245=>"0001001000000011",
                246=>"0001010011111100", 
                247=>"0001100010100000",
                248=>"0001111010111100",
                249=>"0010100001100000",
                250=>"0010001110000011",
                others=>(others=>'0')
                );
begin
   dat<=dato(to_integer(unsigned(add)));
end architecture beh;
